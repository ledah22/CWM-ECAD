//////////////////////////////////////////////////////////////////////////////////
// Exercise #7
// Student Name:ISIDORA RADENKOVIC
// Date: June 5th, 2020
//
//  Description: In this exercise, you need to implement a times table of 0..7x0..7
//  using a memory.
//
//  inputs:
//           clk, a[2:0], b[2:0], read
//
//  outputs:
//           result[4:0]
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns/100ps
module Multiply(
input clk,
input reg [2:0] a,
input reg [2:0] b,
input read,
output reg [4:0] result);


endmodule
